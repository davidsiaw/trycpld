module top (input [1:0]A, output [1:0]Q);
  assign Q = A;
endmodule
