module top (input A, output Q);
  assign Q = A;
endmodule
