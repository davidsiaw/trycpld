module top (input A, output Q);
  INV nn(.A(A), .QN(Q));
endmodule
