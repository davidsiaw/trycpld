module top (input [15:0]A, output [15:0]Q);
  assign Q = A;
endmodule
