module top (input A, output Q);
  INBUF nn(.A(A), .Q(Q));
endmodule
